library verilog;
use verilog.vl_types.all;
entity l2array_sv_unit is
end l2array_sv_unit;
