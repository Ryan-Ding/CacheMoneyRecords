library verilog;
use verilog.vl_types.all;
entity srmask_sv_unit is
end srmask_sv_unit;
