library verilog;
use verilog.vl_types.all;
entity local_br_predictor_sv_unit is
end local_br_predictor_sv_unit;
