library verilog;
use verilog.vl_types.all;
entity br_ctrl_sv_unit is
end br_ctrl_sv_unit;
