library verilog;
use verilog.vl_types.all;
entity add_sv_unit is
end add_sv_unit;
