library verilog;
use verilog.vl_types.all;
entity datapath is
end datapath;
