library verilog;
use verilog.vl_types.all;
entity incremental_counter_sv_unit is
end incremental_counter_sv_unit;
