library verilog;
use verilog.vl_types.all;
entity ewb is
end ewb;
