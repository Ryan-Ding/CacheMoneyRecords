library verilog;
use verilog.vl_types.all;
entity btb_datapath_sv_unit is
end btb_datapath_sv_unit;
