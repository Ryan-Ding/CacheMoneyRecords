library verilog;
use verilog.vl_types.all;
entity global_br_predictor_sv_unit is
end global_br_predictor_sv_unit;
