library verilog;
use verilog.vl_types.all;
entity mem_enable_ctrl_sv_unit is
end mem_enable_ctrl_sv_unit;
