library verilog;
use verilog.vl_types.all;
entity ldi_sti_control_sv_unit is
end ldi_sti_control_sv_unit;
