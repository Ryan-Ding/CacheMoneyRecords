library verilog;
use verilog.vl_types.all;
entity cache_interconnect_datapath_sv_unit is
end cache_interconnect_datapath_sv_unit;
