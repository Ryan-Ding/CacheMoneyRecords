library verilog;
use verilog.vl_types.all;
entity btb_array_sv_unit is
end btb_array_sv_unit;
