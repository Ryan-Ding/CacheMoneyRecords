library verilog;
use verilog.vl_types.all;
entity cache_interconnect is
end cache_interconnect;
