library verilog;
use verilog.vl_types.all;
entity pht_update_ctrl_sv_unit is
end pht_update_ctrl_sv_unit;
