library verilog;
use verilog.vl_types.all;
entity cpudatainmux_sv_unit is
end cpudatainmux_sv_unit;
