library verilog;
use verilog.vl_types.all;
entity \branch_detection__sv_unit\ is
end \branch_detection__sv_unit\;
