library verilog;
use verilog.vl_types.all;
entity mdrmask_sv_unit is
end mdrmask_sv_unit;
