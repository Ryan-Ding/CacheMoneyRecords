library verilog;
use verilog.vl_types.all;
entity choice_predictor_sv_unit is
end choice_predictor_sv_unit;
